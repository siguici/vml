module vml

pub type Translations = map[string]string
pub type GlobalTranslations = map[string]Translations
