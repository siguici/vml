module vml

const entities = [
	'Á',
	'&Aacute;',
	'á',
	'&aacute;',
	'Ă',
	'&Abreve;',
	'ă',
	'&abreve;',
	'∾',
	'&ac;',
	'∿',
	'&acd;',
	'∾̳',
	'&acE;',
	'Â',
	'&Acirc;',
	'â',
	'&acirc;',
	'´',
	'&acute;',
	'А',
	'&Acy;',
	'а',
	'&acy;',
	'Æ',
	'&AElig;',
	'æ',
	'&aelig;',
	'⁡',
	'&af;',
	'𝔄',
	'&Afr;',
	'𝔞',
	'&afr;',
	'À',
	'&Agrave;',
	'à',
	'&agrave;',
	'ℵ',
	'&alefsym;',
	'ℵ',
	'&aleph;',
	'Α',
	'&Alpha;',
	'α',
	'&alpha;',
	'Ā',
	'&Amacr;',
	'ā',
	'&amacr;',
	'⨿',
	'&amalg;',
	'&',
	'&AMP;',
	'&',
	'&amp;',
	'⩓',
	'&And;',
	'∧',
	'&and;',
	'⩕',
	'&andand;',
	'⩜',
	'&andd;',
	'⩘',
	'&andslope;',
	'⩚',
	'&andv;',
	'∠',
	'&ang;',
	'⦤',
	'&ange;',
	'∠',
	'&angle;',
	'∡',
	'&angmsd;',
	'⦨',
	'&angmsdaa;',
	'⦩',
	'&angmsdab;',
	'⦪',
	'&angmsdac;',
	'⦫',
	'&angmsdad;',
	'⦬',
	'&angmsdae;',
	'⦭',
	'&angmsdaf;',
	'⦮',
	'&angmsdag;',
	'⦯',
	'&angmsdah;',
	'∟',
	'&angrt;',
	'⊾',
	'&angrtvb;',
	'⦝',
	'&angrtvbd;',
	'∢',
	'&angsph;',
	'Å',
	'&angst;',
	'⍼',
	'&angzarr;',
	'Ą',
	'&Aogon;',
	'ą',
	'&aogon;',
	'𝔸',
	'&Aopf;',
	'𝕒',
	'&aopf;',
	'≈',
	'&ap;',
	'⩯',
	'&apacir;',
	'⩰',
	'&apE;',
	'≊',
	'&ape;',
	'≋',
	'&apid;',
	"'",
	'&apos;',
	'⁡',
	'&ApplyFunction;',
	'≈',
	'&approx;',
	'≊',
	'&approxeq;',
	'Å',
	'&Aring;',
	'å',
	'&aring;',
	'𝒜',
	'&Ascr;',
	'𝒶',
	'&ascr;',
	'≔',
	'&Assign;',
	'*',
	'&ast;',
	'≈',
	'&asymp;',
	'≍',
	'&asympeq;',
	'Ã',
	'&Atilde;',
	'ã',
	'&atilde;',
	'Ä',
	'&Auml;',
	'ä',
	'&auml;',
	'∳',
	'&awconint;',
	'⨑',
	'&awint;',
	'≌',
	'&backcong;',
	'϶',
	'&backepsilon;',
	'‵',
	'&backprime;',
	'∽',
	'&backsim;',
	'⋍',
	'&backsimeq;',
	'∖',
	'&Backslash;',
	'⫧',
	'&Barv;',
	'⊽',
	'&barvee;',
	'⌆',
	'&Barwed;',
	'⌅',
	'&barwed;',
	'⌅',
	'&barwedge;',
	'⎵',
	'&bbrk;',
	'⎶',
	'&bbrktbrk;',
	'≌',
	'&bcong;',
	'Б',
	'&Bcy;',
	'б',
	'&bcy;',
	'„',
	'&bdquo;',
	'∵',
	'&becaus;',
	'∵',
	'&Because;',
	'∵',
	'&because;',
	'⦰',
	'&bemptyv;',
	'϶',
	'&bepsi;',
	'ℬ',
	'&bernou;',
	'ℬ',
	'&Bernoullis;',
	'Β',
	'&Beta;',
	'β',
	'&beta;',
	'ℶ',
	'&beth;',
	'≬',
	'&between;',
	'𝔅',
	'&Bfr;',
	'𝔟',
	'&bfr;',
	'⋂',
	'&bigcap;',
	'◯',
	'&bigcirc;',
	'⋃',
	'&bigcup;',
	'⨀',
	'&bigodot;',
	'⨁',
	'&bigoplus;',
	'⨂',
	'&bigotimes;',
	'⨆',
	'&bigsqcup;',
	'★',
	'&bigstar;',
	'▽',
	'&bigtriangledown;',
	'△',
	'&bigtriangleup;',
	'⨄',
	'&biguplus;',
	'⋁',
	'&bigvee;',
	'⋀',
	'&bigwedge;',
	'⤍',
	'&bkarow;',
	'⧫',
	'&blacklozenge;',
	'▪',
	'&blacksquare;',
	'▴',
	'&blacktriangle;',
	'▾',
	'&blacktriangledown;',
	'◂',
	'&blacktriangleleft;',
	'▸',
	'&blacktriangleright;',
	'␣',
	'&blank;',
	'▒',
	'&blk12;',
	'░',
	'&blk14;',
	'▓',
	'&blk34;',
	'█',
	'&block;',
	'=⃥',
	'&bne;',
	'≡⃥',
	'&bnequiv;',
	'⫭',
	'&bNot;',
	'⌐',
	'&bnot;',
	'𝔹',
	'&Bopf;',
	'𝕓',
	'&bopf;',
	'⊥',
	'&bot;',
	'⊥',
	'&bottom;',
	'⋈',
	'&bowtie;',
	'⧉',
	'&boxbox;',
	'╗',
	'&boxDL;',
	'╖',
	'&boxDl;',
	'╕',
	'&boxdL;',
	'┐',
	'&boxdl;',
	'╔',
	'&boxDR;',
	'╓',
	'&boxDr;',
	'╒',
	'&boxdR;',
	'┌',
	'&boxdr;',
	'═',
	'&boxH;',
	'─',
	'&boxh;',
	'╦',
	'&boxHD;',
	'╤',
	'&boxHd;',
	'╥',
	'&boxhD;',
	'┬',
	'&boxhd;',
	'╩',
	'&boxHU;',
	'╧',
	'&boxHu;',
	'╨',
	'&boxhU;',
	'┴',
	'&boxhu;',
	'⊟',
	'&boxminus;',
	'⊞',
	'&boxplus;',
	'⊠',
	'&boxtimes;',
	'╝',
	'&boxUL;',
	'╜',
	'&boxUl;',
	'╛',
	'&boxuL;',
	'┘',
	'&boxul;',
	'╚',
	'&boxUR;',
	'╙',
	'&boxUr;',
	'╘',
	'&boxuR;',
	'└',
	'&boxur;',
	'║',
	'&boxV;',
	'│',
	'&boxv;',
	'╬',
	'&boxVH;',
	'╫',
	'&boxVh;',
	'╪',
	'&boxvH;',
	'┼',
	'&boxvh;',
	'╣',
	'&boxVL;',
	'╢',
	'&boxVl;',
	'╡',
	'&boxvL;',
	'┤',
	'&boxvl;',
	'╠',
	'&boxVR;',
	'╟',
	'&boxVr;',
	'╞',
	'&boxvR;',
	'├',
	'&boxvr;',
	'‵',
	'&bprime;',
	'˘',
	'&Breve;',
	'˘',
	'&breve;',
	'¦',
	'&brvbar;',
	'ℬ',
	'&Bscr;',
	'𝒷',
	'&bscr;',
	'⁏',
	'&bsemi;',
	'∽',
	'&bsim;',
	'⋍',
	'&bsime;',
	'\\',
	'&bsol;',
	'⧅',
	'&bsolb;',
	'⟈',
	'&bsolhsub;',
	'•',
	'&bull;',
	'•',
	'&bullet;',
	'≎',
	'&bump;',
	'⪮',
	'&bumpE;',
	'≏',
	'&bumpe;',
	'≎',
	'&Bumpeq;',
	'≏',
	'&bumpeq;',
	'Ć',
	'&Cacute;',
	'ć',
	'&cacute;',
	'⋒',
	'&Cap;',
	'∩',
	'&cap;',
	'⩄',
	'&capand;',
	'⩉',
	'&capbrcup;',
	'⩋',
	'&capcap;',
	'⩇',
	'&capcup;',
	'⩀',
	'&capdot;',
	'ⅅ',
	'&CapitalDifferentialD;',
	'∩︀',
	'&caps;',
	'⁁',
	'&caret;',
	'ˇ',
	'&caron;',
	'ℭ',
	'&Cayleys;',
	'⩍',
	'&ccaps;',
	'Č',
	'&Ccaron;',
	'č',
	'&ccaron;',
	'Ç',
	'&Ccedil;',
	'ç',
	'&ccedil;',
	'Ĉ',
	'&Ccirc;',
	'ĉ',
	'&ccirc;',
	'∰',
	'&Cconint;',
	'⩌',
	'&ccups;',
	'⩐',
	'&ccupssm;',
	'Ċ',
	'&Cdot;',
	'ċ',
	'&cdot;',
	'¸',
	'&cedil;',
	'¸',
	'&Cedilla;',
	'⦲',
	'&cemptyv;',
	'¢',
	'&cent;',
	'·',
	'&CenterDot;',
	'·',
	'&centerdot;',
	'ℭ',
	'&Cfr;',
	'𝔠',
	'&cfr;',
	'Ч',
	'&CHcy;',
	'ч',
	'&chcy;',
	'✓',
	'&check;',
	'✓',
	'&checkmark;',
	'Χ',
	'&Chi;',
	'χ',
	'&chi;',
	'○',
	'&cir;',
	'ˆ',
	'&circ;',
	'≗',
	'&circeq;',
	'↺',
	'&circlearrowleft;',
	'↻',
	'&circlearrowright;',
	'⊛',
	'&circledast;',
	'⊚',
	'&circledcirc;',
	'⊝',
	'&circleddash;',
	'⊙',
	'&CircleDot;',
	'®',
	'&circledR;',
	'Ⓢ',
	'&circledS;',
	'⊖',
	'&CircleMinus;',
	'⊕',
	'&CirclePlus;',
	'⊗',
	'&CircleTimes;',
	'⧃',
	'&cirE;',
	'≗',
	'&cire;',
	'⨐',
	'&cirfnint;',
	'⫯',
	'&cirmid;',
	'⧂',
	'&cirscir;',
	'∲',
	'&ClockwiseContourIntegral;',
	'”',
	'&CloseCurlyDoubleQuote;',
	'’',
	'&CloseCurlyQuote;',
	'♣',
	'&clubs;',
	'♣',
	'&clubsuit;',
	'∷',
	'&Colon;',
	':',
	'&colon;',
	'⩴',
	'&Colone;',
	'≔',
	'&colone;',
	'≔',
	'&coloneq;',
	',',
	'&comma;',
	'@',
	'&commat;',
	'∁',
	'&comp;',
	'∘',
	'&compfn;',
	'∁',
	'&complement;',
	'ℂ',
	'&complexes;',
	'≅',
	'&cong;',
	'⩭',
	'&congdot;',
	'≡',
	'&Congruent;',
	'∯',
	'&Conint;',
	'∮',
	'&conint;',
	'∮',
	'&ContourIntegral;',
	'ℂ',
	'&Copf;',
	'𝕔',
	'&copf;',
	'∐',
	'&coprod;',
	'∐',
	'&Coproduct;',
	'©',
	'&COPY;',
	'©',
	'&copy;',
	'℗',
	'&copysr;',
	'∳',
	'&CounterClockwiseContourIntegral;',
	'↵',
	'&crarr;',
	'⨯',
	'&Cross;',
	'✗',
	'&cross;',
	'𝒞',
	'&Cscr;',
	'𝒸',
	'&cscr;',
	'⫏',
	'&csub;',
	'⫑',
	'&csube;',
	'⫐',
	'&csup;',
	'⫒',
	'&csupe;',
	'⋯',
	'&ctdot;',
	'⤸',
	'&cudarrl;',
	'⤵',
	'&cudarrr;',
	'⋞',
	'&cuepr;',
	'⋟',
	'&cuesc;',
	'↶',
	'&cularr;',
	'⤽',
	'&cularrp;',
	'⋓',
	'&Cup;',
	'∪',
	'&cup;',
	'⩈',
	'&cupbrcap;',
	'≍',
	'&CupCap;',
	'⩆',
	'&cupcap;',
	'⩊',
	'&cupcup;',
	'⊍',
	'&cupdot;',
	'⩅',
	'&cupor;',
	'∪︀',
	'&cups;',
	'↷',
	'&curarr;',
	'⤼',
	'&curarrm;',
	'⋞',
	'&curlyeqprec;',
	'⋟',
	'&curlyeqsucc;',
	'⋎',
	'&curlyvee;',
	'⋏',
	'&curlywedge;',
	'¤',
	'&curren;',
	'↶',
	'&curvearrowleft;',
	'↷',
	'&curvearrowright;',
	'⋎',
	'&cuvee;',
	'⋏',
	'&cuwed;',
	'∲',
	'&cwconint;',
	'∱',
	'&cwint;',
	'⌭',
	'&cylcty;',
	'‡',
	'&Dagger;',
	'†',
	'&dagger;',
	'ℸ',
	'&daleth;',
	'↡',
	'&Darr;',
	'⇓',
	'&dArr;',
	'↓',
	'&darr;',
	'‐',
	'&dash;',
	'⫤',
	'&Dashv;',
	'⊣',
	'&dashv;',
	'⤏',
	'&dbkarow;',
	'˝',
	'&dblac;',
	'Ď',
	'&Dcaron;',
	'ď',
	'&dcaron;',
	'Д',
	'&Dcy;',
	'д',
	'&dcy;',
	'ⅅ',
	'&DD;',
	'ⅆ',
	'&dd;',
	'‡',
	'&ddagger;',
	'⇊',
	'&ddarr;',
	'⤑',
	'&DDotrahd;',
	'⩷',
	'&ddotseq;',
	'°',
	'&deg;',
	'∇',
	'&Del;',
	'Δ',
	'&Delta;',
	'δ',
	'&delta;',
	'⦱',
	'&demptyv;',
	'⥿',
	'&dfisht;',
	'𝔇',
	'&Dfr;',
	'𝔡',
	'&dfr;',
	'⥥',
	'&dHar;',
	'⇃',
	'&dharl;',
	'⇂',
	'&dharr;',
	'´',
	'&DiacriticalAcute;',
	'˙',
	'&DiacriticalDot;',
	'˝',
	'&DiacriticalDoubleAcute;',
	'`',
	'&DiacriticalGrave;',
	'˜',
	'&DiacriticalTilde;',
	'⋄',
	'&diam;',
	'⋄',
	'&Diamond;',
	'⋄',
	'&diamond;',
	'♦',
	'&diamondsuit;',
	'♦',
	'&diams;',
	'¨',
	'&die;',
	'ⅆ',
	'&DifferentialD;',
	'ϝ',
	'&digamma;',
	'⋲',
	'&disin;',
	'÷',
	'&div;',
	'÷',
	'&divide;',
	'⋇',
	'&divideontimes;',
	'⋇',
	'&divonx;',
	'Ђ',
	'&DJcy;',
	'ђ',
	'&djcy;',
	'⌞',
	'&dlcorn;',
	'⌍',
	'&dlcrop;',
	'$',
	'&dollar;',
	'𝔻',
	'&Dopf;',
	'𝕕',
	'&dopf;',
	'¨',
	'&Dot;',
	'˙',
	'&dot;',
	'◌⃜',
	'&DotDot;',
	'≐',
	'&doteq;',
	'≑',
	'&doteqdot;',
	'≐',
	'&DotEqual;',
	'∸',
	'&dotminus;',
	'∔',
	'&dotplus;',
	'⊡',
	'&dotsquare;',
	'⌆',
	'&doublebarwedge;',
	'∯',
	'&DoubleContourIntegral;',
	'¨',
	'&DoubleDot;',
	'⇓',
	'&DoubleDownArrow;',
	'⇐',
	'&DoubleLeftArrow;',
	'⇔',
	'&DoubleLeftRightArrow;',
	'⫤',
	'&DoubleLeftTee;',
	'⟸',
	'&DoubleLongLeftArrow;',
	'⟺',
	'&DoubleLongLeftRightArrow;',
	'⟹',
	'&DoubleLongRightArrow;',
	'⇒',
	'&DoubleRightArrow;',
	'⊨',
	'&DoubleRightTee;',
	'⇑',
	'&DoubleUpArrow;',
	'⇕',
	'&DoubleUpDownArrow;',
	'∥',
	'&DoubleVerticalBar;',
	'↓',
	'&DownArrow;',
	'⇓',
	'&Downarrow;',
	'↓',
	'&downarrow;',
	'⤓',
	'&DownArrowBar;',
	'⇵',
	'&DownArrowUpArrow;',
	'◌̑',
	'&DownBreve;',
	'⇊',
	'&downdownarrows;',
	'⇃',
	'&downharpoonleft;',
	'⇂',
	'&downharpoonright;',
	'⥐',
	'&DownLeftRightVector;',
	'⥞',
	'&DownLeftTeeVector;',
	'↽',
	'&DownLeftVector;',
	'⥖',
	'&DownLeftVectorBar;',
	'⥟',
	'&DownRightTeeVector;',
	'⇁',
	'&DownRightVector;',
	'⥗',
	'&DownRightVectorBar;',
	'⊤',
	'&DownTee;',
	'↧',
	'&DownTeeArrow;',
	'⤐',
	'&drbkarow;',
	'⌟',
	'&drcorn;',
	'⌌',
	'&drcrop;',
	'𝒟',
	'&Dscr;',
	'𝒹',
	'&dscr;',
	'Ѕ',
	'&DScy;',
	'ѕ',
	'&dscy;',
	'⧶',
	'&dsol;',
	'Đ',
	'&Dstrok;',
	'đ',
	'&dstrok;',
	'⋱',
	'&dtdot;',
	'▿',
	'&dtri;',
	'▾',
	'&dtrif;',
	'⇵',
	'&duarr;',
	'⥯',
	'&duhar;',
	'⦦',
	'&dwangle;',
	'Џ',
	'&DZcy;',
	'џ',
	'&dzcy;',
	'⟿',
	'&dzigrarr;',
	'É',
	'&Eacute;',
	'é',
	'&eacute;',
	'⩮',
	'&easter;',
	'Ě',
	'&Ecaron;',
	'ě',
	'&ecaron;',
	'≖',
	'&ecir;',
	'Ê',
	'&Ecirc;',
	'ê',
	'&ecirc;',
	'≕',
	'&ecolon;',
	'Э',
	'&Ecy;',
	'э',
	'&ecy;',
	'⩷',
	'&eDDot;',
	'Ė',
	'&Edot;',
	'≑',
	'&eDot;',
	'ė',
	'&edot;',
	'ⅇ',
	'&ee;',
	'≒',
	'&efDot;',
	'𝔈',
	'&Efr;',
	'𝔢',
	'&efr;',
	'⪚',
	'&eg;',
	'È',
	'&Egrave;',
	'è',
	'&egrave;',
	'⪖',
	'&egs;',
	'⪘',
	'&egsdot;',
	'⪙',
	'&el;',
	'∈',
	'&Element;',
	'⏧',
	'&elinters;',
	'ℓ',
	'&ell;',
	'⪕',
	'&els;',
	'⪗',
	'&elsdot;',
	'Ē',
	'&Emacr;',
	'ē',
	'&emacr;',
	'∅',
	'&empty;',
	'∅',
	'&emptyset;',
	'◻',
	'&EmptySmallSquare;',
	'∅',
	'&emptyv;',
	'▫',
	'&EmptyVerySmallSquare;',
	' ',
	'&emsp;',
	' ',
	'&emsp13;',
	' ',
	'&emsp14;',
	'Ŋ',
	'&ENG;',
	'ŋ',
	'&eng;',
	' ',
	'&ensp;',
	'Ę',
	'&Eogon;',
	'ę',
	'&eogon;',
	'𝔼',
	'&Eopf;',
	'𝕖',
	'&eopf;',
	'⋕',
	'&epar;',
	'⧣',
	'&eparsl;',
	'⩱',
	'&eplus;',
	'ε',
	'&epsi;',
	'Ε',
	'&Epsilon;',
	'ε',
	'&epsilon;',
	'ϵ',
	'&epsiv;',
	'≖',
	'&eqcirc;',
	'≕',
	'&eqcolon;',
	'≂',
	'&eqsim;',
	'⪖',
	'&eqslantgtr;',
	'⪕',
	'&eqslantless;',
	'⩵',
	'&Equal;',
	'=',
	'&equals;',
	'≂',
	'&EqualTilde;',
	'≟',
	'&equest;',
	'⇌',
	'&Equilibrium;',
	'≡',
	'&equiv;',
	'⩸',
	'&equivDD;',
	'⧥',
	'&eqvparsl;',
	'⥱',
	'&erarr;',
	'≓',
	'&erDot;',
	'ℰ',
	'&Escr;',
	'ℯ',
	'&escr;',
	'≐',
	'&esdot;',
	'⩳',
	'&Esim;',
	'≂',
	'&esim;',
	'Η',
	'&Eta;',
	'η',
	'&eta;',
	'Ð',
	'&ETH;',
	'ð',
	'&eth;',
	'Ë',
	'&Euml;',
	'ë',
	'&euml;',
	'€',
	'&euro;',
	'!',
	'&excl;',
	'∃',
	'&exist;',
	'∃',
	'&Exists;',
	'ℰ',
	'&expectation;',
	'ⅇ',
	'&ExponentialE;',
	'ⅇ',
	'&exponentiale;',
	'≒',
	'&fallingdotseq;',
	'Ф',
	'&Fcy;',
	'ф',
	'&fcy;',
	'♀',
	'&female;',
	'ﬃ',
	'&ffilig;',
	'ﬀ',
	'&fflig;',
	'ﬄ',
	'&ffllig;',
	'𝔉',
	'&Ffr;',
	'𝔣',
	'&ffr;',
	'ﬁ',
	'&filig;',
	'◼',
	'&FilledSmallSquare;',
	'▪',
	'&FilledVerySmallSquare;',
	'fj',
	'&fjlig;',
	'♭',
	'&flat;',
	'ﬂ',
	'&fllig;',
	'▱',
	'&fltns;',
	'ƒ',
	'&fnof;',
	'𝔽',
	'&Fopf;',
	'𝕗',
	'&fopf;',
	'∀',
	'&ForAll;',
	'∀',
	'&forall;',
	'⋔',
	'&fork;',
	'⫙',
	'&forkv;',
	'ℱ',
	'&Fouriertrf;',
	'⨍',
	'&fpartint;',
	'½',
	'&frac12;',
	'⅓',
	'&frac13;',
	'¼',
	'&frac14;',
	'⅕',
	'&frac15;',
	'⅙',
	'&frac16;',
	'⅛',
	'&frac18;',
	'⅔',
	'&frac23;',
	'⅖',
	'&frac25;',
	'¾',
	'&frac34;',
	'⅗',
	'&frac35;',
	'⅜',
	'&frac38;',
	'⅘',
	'&frac45;',
	'⅚',
	'&frac56;',
	'⅝',
	'&frac58;',
	'⅞',
	'&frac78;',
	'⁄',
	'&frasl;',
	'⌢',
	'&frown;',
	'ℱ',
	'&Fscr;',
	'𝒻',
	'&fscr;',
	'ǵ',
	'&gacute;',
	'Γ',
	'&Gamma;',
	'γ',
	'&gamma;',
	'Ϝ',
	'&Gammad;',
	'ϝ',
	'&gammad;',
	'⪆',
	'&gap;',
	'Ğ',
	'&Gbreve;',
	'ğ',
	'&gbreve;',
	'Ģ',
	'&Gcedil;',
	'Ĝ',
	'&Gcirc;',
	'ĝ',
	'&gcirc;',
	'Г',
	'&Gcy;',
	'г',
	'&gcy;',
	'Ġ',
	'&Gdot;',
	'ġ',
	'&gdot;',
	'≧',
	'&gE;',
	'≥',
	'&ge;',
	'⪌',
	'&gEl;',
	'⋛',
	'&gel;',
	'≥',
	'&geq;',
	'≧',
	'&geqq;',
	'⩾',
	'&geqslant;',
	'⩾',
	'&ges;',
	'⪩',
	'&gescc;',
	'⪀',
	'&gesdot;',
	'⪂',
	'&gesdoto;',
	'⪄',
	'&gesdotol;',
	'⋛︀',
	'&gesl;',
	'⪔',
	'&gesles;',
	'𝔊',
	'&Gfr;',
	'𝔤',
	'&gfr;',
	'⋙',
	'&Gg;',
	'≫',
	'&gg;',
	'⋙',
	'&ggg;',
	'ℷ',
	'&gimel;',
	'Ѓ',
	'&GJcy;',
	'ѓ',
	'&gjcy;',
	'≷',
	'&gl;',
	'⪥',
	'&gla;',
	'⪒',
	'&glE;',
	'⪤',
	'&glj;',
	'⪊',
	'&gnap;',
	'⪊',
	'&gnapprox;',
	'≩',
	'&gnE;',
	'⪈',
	'&gne;',
	'⪈',
	'&gneq;',
	'≩',
	'&gneqq;',
	'⋧',
	'&gnsim;',
	'𝔾',
	'&Gopf;',
	'𝕘',
	'&gopf;',
	'`',
	'&grave;',
	'≥',
	'&GreaterEqual;',
	'⋛',
	'&GreaterEqualLess;',
	'≧',
	'&GreaterFullEqual;',
	'⪢',
	'&GreaterGreater;',
	'≷',
	'&GreaterLess;',
	'⩾',
	'&GreaterSlantEqual;',
	'≳',
	'&GreaterTilde;',
	'𝒢',
	'&Gscr;',
	'ℊ',
	'&gscr;',
	'≳',
	'&gsim;',
	'⪎',
	'&gsime;',
	'⪐',
	'&gsiml;',
	'>',
	'&GT;',
	'≫',
	'&Gt;',
	'>',
	'&gt;',
	'⪧',
	'&gtcc;',
	'⩺',
	'&gtcir;',
	'⋗',
	'&gtdot;',
	'⦕',
	'&gtlPar;',
	'⩼',
	'&gtquest;',
	'⪆',
	'&gtrapprox;',
	'⥸',
	'&gtrarr;',
	'⋗',
	'&gtrdot;',
	'⋛',
	'&gtreqless;',
	'⪌',
	'&gtreqqless;',
	'≷',
	'&gtrless;',
	'≳',
	'&gtrsim;',
	'≩︀',
	'&gvertneqq;',
	'≩︀',
	'&gvnE;',
	'ˇ',
	'&Hacek;',
	' ',
	'&hairsp;',
	'½',
	'&half;',
	'ℋ',
	'&hamilt;',
	'Ъ',
	'&HARDcy;',
	'ъ',
	'&hardcy;',
	'⇔',
	'&hArr;',
	'↔',
	'&harr;',
	'⥈',
	'&harrcir;',
	'↭',
	'&harrw;',
	'^',
	'&Hat;',
	'ℏ',
	'&hbar;',
	'Ĥ',
	'&Hcirc;',
	'ĥ',
	'&hcirc;',
	'♥',
	'&hearts;',
	'♥',
	'&heartsuit;',
	'…',
	'&hellip;',
	'⊹',
	'&hercon;',
	'ℌ',
	'&Hfr;',
	'𝔥',
	'&hfr;',
	'ℋ',
	'&HilbertSpace;',
	'⤥',
	'&hksearow;',
	'⤦',
	'&hkswarow;',
	'⇿',
	'&hoarr;',
	'∻',
	'&homtht;',
	'↩',
	'&hookleftarrow;',
	'↪',
	'&hookrightarrow;',
	'ℍ',
	'&Hopf;',
	'𝕙',
	'&hopf;',
	'―',
	'&horbar;',
	'─',
	'&HorizontalLine;',
	'ℋ',
	'&Hscr;',
	'𝒽',
	'&hscr;',
	'ℏ',
	'&hslash;',
	'Ħ',
	'&Hstrok;',
	'ħ',
	'&hstrok;',
	'≎',
	'&HumpDownHump;',
	'≏',
	'&HumpEqual;',
	'⁃',
	'&hybull;',
	'‐',
	'&hyphen;',
	'Í',
	'&Iacute;',
	'í',
	'&iacute;',
	'⁣',
	'&ic;',
	'Î',
	'&Icirc;',
	'î',
	'&icirc;',
	'И',
	'&Icy;',
	'и',
	'&icy;',
	'İ',
	'&Idot;',
	'Е',
	'&IEcy;',
	'е',
	'&iecy;',
	'¡',
	'&iexcl;',
	'⇔',
	'&iff;',
	'ℑ',
	'&Ifr;',
	'𝔦',
	'&ifr;',
	'Ì',
	'&Igrave;',
	'ì',
	'&igrave;',
	'ⅈ',
	'&ii;',
	'⨌',
	'&iiiint;',
	'∭',
	'&iiint;',
	'⧜',
	'&iinfin;',
	'℩',
	'&iiota;',
	'Ĳ',
	'&IJlig;',
	'ĳ',
	'&ijlig;',
	'ℑ',
	'&Im;',
	'Ī',
	'&Imacr;',
	'ī',
	'&imacr;',
	'ℑ',
	'&image;',
	'ⅈ',
	'&ImaginaryI;',
	'ℐ',
	'&imagline;',
	'ℑ',
	'&imagpart;',
	'ı',
	'&imath;',
	'⊷',
	'&imof;',
	'Ƶ',
	'&imped;',
	'⇒',
	'&Implies;',
	'∈',
	'&in;',
	'℅',
	'&incare;',
	'∞',
	'&infin;',
	'⧝',
	'&infintie;',
	'ı',
	'&inodot;',
	'∬',
	'&Int;',
	'∫',
	'&int;',
	'⊺',
	'&intcal;',
	'ℤ',
	'&integers;',
	'∫',
	'&Integral;',
	'⊺',
	'&intercal;',
	'⋂',
	'&Intersection;',
	'⨗',
	'&intlarhk;',
	'⨼',
	'&intprod;',
	'⁣',
	'&InvisibleComma;',
	'⁢',
	'&InvisibleTimes;',
	'Ё',
	'&IOcy;',
	'ё',
	'&iocy;',
	'Į',
	'&Iogon;',
	'į',
	'&iogon;',
	'𝕀',
	'&Iopf;',
	'𝕚',
	'&iopf;',
	'Ι',
	'&Iota;',
	'ι',
	'&iota;',
	'⨼',
	'&iprod;',
	'¿',
	'&iquest;',
	'ℐ',
	'&Iscr;',
	'𝒾',
	'&iscr;',
	'∈',
	'&isin;',
	'⋵',
	'&isindot;',
	'⋹',
	'&isinE;',
	'⋴',
	'&isins;',
	'⋳',
	'&isinsv;',
	'∈',
	'&isinv;',
	'⁢',
	'&it;',
	'Ĩ',
	'&Itilde;',
	'ĩ',
	'&itilde;',
	'І',
	'&Iukcy;',
	'і',
	'&iukcy;',
	'Ï',
	'&Iuml;',
	'ï',
	'&iuml;',
	'Ĵ',
	'&Jcirc;',
	'ĵ',
	'&jcirc;',
	'Й',
	'&Jcy;',
	'й',
	'&jcy;',
	'𝔍',
	'&Jfr;',
	'𝔧',
	'&jfr;',
	'ȷ',
	'&jmath;',
	'𝕁',
	'&Jopf;',
	'𝕛',
	'&jopf;',
	'𝒥',
	'&Jscr;',
	'𝒿',
	'&jscr;',
	'Ј',
	'&Jsercy;',
	'ј',
	'&jsercy;',
	'Є',
	'&Jukcy;',
	'є',
	'&jukcy;',
	'Κ',
	'&Kappa;',
	'κ',
	'&kappa;',
	'ϰ',
	'&kappav;',
	'Ķ',
	'&Kcedil;',
	'ķ',
	'&kcedil;',
	'К',
	'&Kcy;',
	'к',
	'&kcy;',
	'𝔎',
	'&Kfr;',
	'𝔨',
	'&kfr;',
	'ĸ',
	'&kgreen;',
	'Х',
	'&KHcy;',
	'х',
	'&khcy;',
	'Ќ',
	'&KJcy;',
	'ќ',
	'&kjcy;',
	'𝕂',
	'&Kopf;',
	'𝕜',
	'&kopf;',
	'𝒦',
	'&Kscr;',
	'𝓀',
	'&kscr;',
	'⇚',
	'&lAarr;',
	'Ĺ',
	'&Lacute;',
	'ĺ',
	'&lacute;',
	'⦴',
	'&laemptyv;',
	'ℒ',
	'&lagran;',
	'Λ',
	'&Lambda;',
	'λ',
	'&lambda;',
	'⟪',
	'&Lang;',
	'⟨',
	'&lang;',
	'⦑',
	'&langd;',
	'⟨',
	'&langle;',
	'⪅',
	'&lap;',
	'ℒ',
	'&Laplacetrf;',
	'«',
	'&laquo;',
	'↞',
	'&Larr;',
	'⇐',
	'&lArr;',
	'←',
	'&larr;',
	'⇤',
	'&larrb;',
	'⤟',
	'&larrbfs;',
	'⤝',
	'&larrfs;',
	'↩',
	'&larrhk;',
	'↫',
	'&larrlp;',
	'⤹',
	'&larrpl;',
	'⥳',
	'&larrsim;',
	'↢',
	'&larrtl;',
	'⪫',
	'&lat;',
	'⤛',
	'&lAtail;',
	'⤙',
	'&latail;',
	'⪭',
	'&late;',
	'⪭︀',
	'&lates;',
	'⤎',
	'&lBarr;',
	'⤌',
	'&lbarr;',
	'❲',
	'&lbbrk;',
	'{',
	'&lbrace;',
	'[',
	'&lbrack;',
	'⦋',
	'&lbrke;',
	'⦏',
	'&lbrksld;',
	'⦍',
	'&lbrkslu;',
	'Ľ',
	'&Lcaron;',
	'ľ',
	'&lcaron;',
	'Ļ',
	'&Lcedil;',
	'ļ',
	'&lcedil;',
	'⌈',
	'&lceil;',
	'{',
	'&lcub;',
	'Л',
	'&Lcy;',
	'л',
	'&lcy;',
	'⤶',
	'&ldca;',
	'“',
	'&ldquo;',
	'„',
	'&ldquor;',
	'⥧',
	'&ldrdhar;',
	'⥋',
	'&ldrushar;',
	'↲',
	'&ldsh;',
	'≦',
	'&lE;',
	'≤',
	'&le;',
	'⟨',
	'&LeftAngleBracket;',
	'←',
	'&LeftArrow;',
	'⇐',
	'&Leftarrow;',
	'←',
	'&leftarrow;',
	'⇤',
	'&LeftArrowBar;',
	'⇆',
	'&LeftArrowRightArrow;',
	'↢',
	'&leftarrowtail;',
	'⌈',
	'&LeftCeiling;',
	'⟦',
	'&LeftDoubleBracket;',
	'⥡',
	'&LeftDownTeeVector;',
	'⇃',
	'&LeftDownVector;',
	'⥙',
	'&LeftDownVectorBar;',
	'⌊',
	'&LeftFloor;',
	'↽',
	'&leftharpoondown;',
	'↼',
	'&leftharpoonup;',
	'⇇',
	'&leftleftarrows;',
	'↔',
	'&LeftRightArrow;',
	'⇔',
	'&Leftrightarrow;',
	'↔',
	'&leftrightarrow;',
	'⇆',
	'&leftrightarrows;',
	'⇋',
	'&leftrightharpoons;',
	'↭',
	'&leftrightsquigarrow;',
	'⥎',
	'&LeftRightVector;',
	'⊣',
	'&LeftTee;',
	'↤',
	'&LeftTeeArrow;',
	'⥚',
	'&LeftTeeVector;',
	'⋋',
	'&leftthreetimes;',
	'⊲',
	'&LeftTriangle;',
	'⧏',
	'&LeftTriangleBar;',
	'⊴',
	'&LeftTriangleEqual;',
	'⥑',
	'&LeftUpDownVector;',
	'⥠',
	'&LeftUpTeeVector;',
	'↿',
	'&LeftUpVector;',
	'⥘',
	'&LeftUpVectorBar;',
	'↼',
	'&LeftVector;',
	'⥒',
	'&LeftVectorBar;',
	'⪋',
	'&lEg;',
	'⋚',
	'&leg;',
	'≤',
	'&leq;',
	'≦',
	'&leqq;',
	'⩽',
	'&leqslant;',
	'⩽',
	'&les;',
	'⪨',
	'&lescc;',
	'⩿',
	'&lesdot;',
	'⪁',
	'&lesdoto;',
	'⪃',
	'&lesdotor;',
	'⋚︀',
	'&lesg;',
	'⪓',
	'&lesges;',
	'⪅',
	'&lessapprox;',
	'⋖',
	'&lessdot;',
	'⋚',
	'&lesseqgtr;',
	'⪋',
	'&lesseqqgtr;',
	'⋚',
	'&LessEqualGreater;',
	'≦',
	'&LessFullEqual;',
	'≶',
	'&LessGreater;',
	'≶',
	'&lessgtr;',
	'⪡',
	'&LessLess;',
	'≲',
	'&lesssim;',
	'⩽',
	'&LessSlantEqual;',
	'≲',
	'&LessTilde;',
	'⥼',
	'&lfisht;',
	'⌊',
	'&lfloor;',
	'𝔏',
	'&Lfr;',
	'𝔩',
	'&lfr;',
	'≶',
	'&lg;',
	'⪑',
	'&lgE;',
	'⥢',
	'&lHar;',
	'↽',
	'&lhard;',
	'↼',
	'&lharu;',
	'⥪',
	'&lharul;',
	'▄',
	'&lhblk;',
	'Љ',
	'&LJcy;',
	'љ',
	'&ljcy;',
	'⋘',
	'&Ll;',
	'≪',
	'&ll;',
	'⇇',
	'&llarr;',
	'⌞',
	'&llcorner;',
	'⇚',
	'&Lleftarrow;',
	'⥫',
	'&llhard;',
	'◺',
	'&lltri;',
	'Ŀ',
	'&Lmidot;',
	'ŀ',
	'&lmidot;',
	'⎰',
	'&lmoust;',
	'⎰',
	'&lmoustache;',
	'⪉',
	'&lnap;',
	'⪉',
	'&lnapprox;',
	'≨',
	'&lnE;',
	'⪇',
	'&lne;',
	'⪇',
	'&lneq;',
	'≨',
	'&lneqq;',
	'⋦',
	'&lnsim;',
	'⟬',
	'&loang;',
	'⇽',
	'&loarr;',
	'⟦',
	'&lobrk;',
	'⟵',
	'&LongLeftArrow;',
	'⟸',
	'&Longleftarrow;',
	'⟵',
	'&longleftarrow;',
	'⟷',
	'&LongLeftRightArrow;',
	'⟺',
	'&Longleftrightarrow;',
	'⟷',
	'&longleftrightarrow;',
	'⟼',
	'&longmapsto;',
	'⟶',
	'&LongRightArrow;',
	'⟹',
	'&Longrightarrow;',
	'⟶',
	'&longrightarrow;',
	'↫',
	'&looparrowleft;',
	'↬',
	'&looparrowright;',
	'⦅',
	'&lopar;',
	'𝕃',
	'&Lopf;',
	'𝕝',
	'&lopf;',
	'⨭',
	'&loplus;',
	'⨴',
	'&lotimes;',
	'∗',
	'&lowast;',
	'_',
	'&lowbar;',
	'↙',
	'&LowerLeftArrow;',
	'↘',
	'&LowerRightArrow;',
	'◊',
	'&loz;',
	'◊',
	'&lozenge;',
	'⧫',
	'&lozf;',
	'(',
	'&lpar;',
	'⦓',
	'&lparlt;',
	'⇆',
	'&lrarr;',
	'⌟',
	'&lrcorner;',
	'⇋',
	'&lrhar;',
	'⥭',
	'&lrhard;',
	'‎',
	'&lrm;',
	'⊿',
	'&lrtri;',
	'‹',
	'&lsaquo;',
	'ℒ',
	'&Lscr;',
	'𝓁',
	'&lscr;',
	'↰',
	'&Lsh;',
	'↰',
	'&lsh;',
	'≲',
	'&lsim;',
	'⪍',
	'&lsime;',
	'⪏',
	'&lsimg;',
	'[',
	'&lsqb;',
	'‘',
	'&lsquo;',
	'‚',
	'&lsquor;',
	'Ł',
	'&Lstrok;',
	'ł',
	'&lstrok;',
	'<',
	'&LT;',
	'≪',
	'&Lt;',
	'<',
	'&lt;',
	'⪦',
	'&ltcc;',
	'⩹',
	'&ltcir;',
	'⋖',
	'&ltdot;',
	'⋋',
	'&lthree;',
	'⋉',
	'&ltimes;',
	'⥶',
	'&ltlarr;',
	'⩻',
	'&ltquest;',
	'◃',
	'&ltri;',
	'⊴',
	'&ltrie;',
	'◂',
	'&ltrif;',
	'⦖',
	'&ltrPar;',
	'⥊',
	'&lurdshar;',
	'⥦',
	'&luruhar;',
	'≨︀',
	'&lvertneqq;',
	'≨︀',
	'&lvnE;',
	'¯',
	'&macr;',
	'♂',
	'&male;',
	'✠',
	'&malt;',
	'✠',
	'&maltese;',
	'⤅',
	'&Map;',
	'↦',
	'&map;',
	'↦',
	'&mapsto;',
	'↧',
	'&mapstodown;',
	'↤',
	'&mapstoleft;',
	'↥',
	'&mapstoup;',
	'▮',
	'&marker;',
	'⨩',
	'&mcomma;',
	'М',
	'&Mcy;',
	'м',
	'&mcy;',
	'—',
	'&mdash;',
	'∺',
	'&mDDot;',
	'∡',
	'&measuredangle;',
	' ',
	'&MediumSpace;',
	'ℳ',
	'&Mellintrf;',
	'𝔐',
	'&Mfr;',
	'𝔪',
	'&mfr;',
	'℧',
	'&mho;',
	'µ',
	'&micro;',
	'∣',
	'&mid;',
	'*',
	'&midast;',
	'⫰',
	'&midcir;',
	'·',
	'&middot;',
	'−',
	'&minus;',
	'⊟',
	'&minusb;',
	'∸',
	'&minusd;',
	'⨪',
	'&minusdu;',
	'∓',
	'&MinusPlus;',
	'⫛',
	'&mlcp;',
	'…',
	'&mldr;',
	'∓',
	'&mnplus;',
	'⊧',
	'&models;',
	'𝕄',
	'&Mopf;',
	'𝕞',
	'&mopf;',
	'∓',
	'&mp;',
	'ℳ',
	'&Mscr;',
	'𝓂',
	'&mscr;',
	'∾',
	'&mstpos;',
	'Μ',
	'&Mu;',
	'μ',
	'&mu;',
	'⊸',
	'&multimap;',
	'⊸',
	'&mumap;',
	'∇',
	'&nabla;',
	'Ń',
	'&Nacute;',
	'ń',
	'&nacute;',
	'∠⃒',
	'&nang;',
	'≉',
	'&nap;',
	'⩰̸',
	'&napE;',
	'≋̸',
	'&napid;',
	'ŉ',
	'&napos;',
	'≉',
	'&napprox;',
	'♮',
	'&natur;',
	'♮',
	'&natural;',
	'ℕ',
	'&naturals;',
	' ',
	'&nbsp;',
	'≎̸',
	'&nbump;',
	'≏̸',
	'&nbumpe;',
	'⩃',
	'&ncap;',
	'Ň',
	'&Ncaron;',
	'ň',
	'&ncaron;',
	'Ņ',
	'&Ncedil;',
	'ņ',
	'&ncedil;',
	'≇',
	'&ncong;',
	'⩭̸',
	'&ncongdot;',
	'⩂',
	'&ncup;',
	'Н',
	'&Ncy;',
	'н',
	'&ncy;',
	'–',
	'&ndash;',
	'≠',
	'&ne;',
	'⤤',
	'&nearhk;',
	'⇗',
	'&neArr;',
	'↗',
	'&nearr;',
	'↗',
	'&nearrow;',
	'≐̸',
	'&nedot;',
	'​',
	'&NegativeMediumSpace;',
	'​',
	'&NegativeThickSpace;',
	'​',
	'&NegativeThinSpace;',
	'​',
	'&NegativeVeryThinSpace;',
	'≢',
	'&nequiv;',
	'⤨',
	'&nesear;',
	'≂̸',
	'&nesim;',
	'≫',
	'&NestedGreaterGreater;',
	'≪',
	'&NestedLessLess;',
	'␊',
	'&NewLine;',
	'∄',
	'&nexist;',
	'∄',
	'&nexists;',
	'𝔑',
	'&Nfr;',
	'𝔫',
	'&nfr;',
	'≧̸',
	'&ngE;',
	'≱',
	'&nge;',
	'≱',
	'&ngeq;',
	'≧̸',
	'&ngeqq;',
	'⩾̸',
	'&ngeqslant;',
	'⩾̸',
	'&nges;',
	'⋙̸',
	'&nGg;',
	'≵',
	'&ngsim;',
	'≫⃒',
	'&nGt;',
	'≯',
	'&ngt;',
	'≯',
	'&ngtr;',
	'≫̸',
	'&nGtv;',
	'⇎',
	'&nhArr;',
	'↮',
	'&nharr;',
	'⫲',
	'&nhpar;',
	'∋',
	'&ni;',
	'⋼',
	'&nis;',
	'⋺',
	'&nisd;',
	'∋',
	'&niv;',
	'Њ',
	'&NJcy;',
	'њ',
	'&njcy;',
	'⇍',
	'&nlArr;',
	'↚',
	'&nlarr;',
	'‥',
	'&nldr;',
	'≦̸',
	'&nlE;',
	'≰',
	'&nle;',
	'⇍',
	'&nLeftarrow;',
	'↚',
	'&nleftarrow;',
	'⇎',
	'&nLeftrightarrow;',
	'↮',
	'&nleftrightarrow;',
	'≰',
	'&nleq;',
	'≦̸',
	'&nleqq;',
	'⩽̸',
	'&nleqslant;',
	'⩽̸',
	'&nles;',
	'≮',
	'&nless;',
	'⋘̸',
	'&nLl;',
	'≴',
	'&nlsim;',
	'≪⃒',
	'&nLt;',
	'≮',
	'&nlt;',
	'⋪',
	'&nltri;',
	'⋬',
	'&nltrie;',
	'≪̸',
	'&nLtv;',
	'∤',
	'&nmid;',
	'⁠',
	'&NoBreak;',
	' ',
	'&NonBreakingSpace;',
	'ℕ',
	'&Nopf;',
	'𝕟',
	'&nopf;',
	'⫬',
	'&Not;',
	'¬',
	'&not;',
	'≢',
	'&NotCongruent;',
	'≭',
	'&NotCupCap;',
	'∦',
	'&NotDoubleVerticalBar;',
	'∉',
	'&NotElement;',
	'≠',
	'&NotEqual;',
	'≂̸',
	'&NotEqualTilde;',
	'∄',
	'&NotExists;',
	'≯',
	'&NotGreater;',
	'≱',
	'&NotGreaterEqual;',
	'≧̸',
	'&NotGreaterFullEqual;',
	'≫̸',
	'&NotGreaterGreater;',
	'≹',
	'&NotGreaterLess;',
	'⩾̸',
	'&NotGreaterSlantEqual;',
	'≵',
	'&NotGreaterTilde;',
	'≎̸',
	'&NotHumpDownHump;',
	'≏̸',
	'&NotHumpEqual;',
	'∉',
	'&notin;',
	'⋵̸',
	'&notindot;',
	'⋹̸',
	'&notinE;',
	'∉',
	'&notinva;',
	'⋷',
	'&notinvb;',
	'⋶',
	'&notinvc;',
	'⋪',
	'&NotLeftTriangle;',
	'⧏̸',
	'&NotLeftTriangleBar;',
	'⋬',
	'&NotLeftTriangleEqual;',
	'≮',
	'&NotLess;',
	'≰',
	'&NotLessEqual;',
	'≸',
	'&NotLessGreater;',
	'≪̸',
	'&NotLessLess;',
	'⩽̸',
	'&NotLessSlantEqual;',
	'≴',
	'&NotLessTilde;',
	'⪢̸',
	'&NotNestedGreaterGreater;',
	'⪡̸',
	'&NotNestedLessLess;',
	'∌',
	'&notni;',
	'∌',
	'&notniva;',
	'⋾',
	'&notnivb;',
	'⋽',
	'&notnivc;',
	'⊀',
	'&NotPrecedes;',
	'⪯̸',
	'&NotPrecedesEqual;',
	'⋠',
	'&NotPrecedesSlantEqual;',
	'∌',
	'&NotReverseElement;',
	'⋫',
	'&NotRightTriangle;',
	'⧐̸',
	'&NotRightTriangleBar;',
	'⋭',
	'&NotRightTriangleEqual;',
	'⊏̸',
	'&NotSquareSubset;',
	'⋢',
	'&NotSquareSubsetEqual;',
	'⊐̸',
	'&NotSquareSuperset;',
	'⋣',
	'&NotSquareSupersetEqual;',
	'⊂⃒',
	'&NotSubset;',
	'⊈',
	'&NotSubsetEqual;',
	'⊁',
	'&NotSucceeds;',
	'⪰̸',
	'&NotSucceedsEqual;',
	'⋡',
	'&NotSucceedsSlantEqual;',
	'≿̸',
	'&NotSucceedsTilde;',
	'⊃⃒',
	'&NotSuperset;',
	'⊉',
	'&NotSupersetEqual;',
	'≁',
	'&NotTilde;',
	'≄',
	'&NotTildeEqual;',
	'≇',
	'&NotTildeFullEqual;',
	'≉',
	'&NotTildeTilde;',
	'∤',
	'&NotVerticalBar;',
	'∦',
	'&npar;',
	'∦',
	'&nparallel;',
	'⫽⃥',
	'&nparsl;',
	'∂̸',
	'&npart;',
	'⨔',
	'&npolint;',
	'⊀',
	'&npr;',
	'⋠',
	'&nprcue;',
	'⪯̸',
	'&npre;',
	'⊀',
	'&nprec;',
	'⪯̸',
	'&npreceq;',
	'⇏',
	'&nrArr;',
	'↛',
	'&nrarr;',
	'⤳̸',
	'&nrarrc;',
	'↝̸',
	'&nrarrw;',
	'⇏',
	'&nRightarrow;',
	'↛',
	'&nrightarrow;',
	'⋫',
	'&nrtri;',
	'⋭',
	'&nrtrie;',
	'⊁',
	'&nsc;',
	'⋡',
	'&nsccue;',
	'⪰̸',
	'&nsce;',
	'𝒩',
	'&Nscr;',
	'𝓃',
	'&nscr;',
	'∤',
	'&nshortmid;',
	'∦',
	'&nshortparallel;',
	'≁',
	'&nsim;',
	'≄',
	'&nsime;',
	'≄',
	'&nsimeq;',
	'∤',
	'&nsmid;',
	'∦',
	'&nspar;',
	'⋢',
	'&nsqsube;',
	'⋣',
	'&nsqsupe;',
	'⊄',
	'&nsub;',
	'⫅̸',
	'&nsubE;',
	'⊈',
	'&nsube;',
	'⊂⃒',
	'&nsubset;',
	'⊈',
	'&nsubseteq;',
	'⫅̸',
	'&nsubseteqq;',
	'⊁',
	'&nsucc;',
	'⪰̸',
	'&nsucceq;',
	'⊅',
	'&nsup;',
	'⫆̸',
	'&nsupE;',
	'⊉',
	'&nsupe;',
	'⊃⃒',
	'&nsupset;',
	'⊉',
	'&nsupseteq;',
	'⫆̸',
	'&nsupseteqq;',
	'≹',
	'&ntgl;',
	'Ñ',
	'&Ntilde;',
	'ñ',
	'&ntilde;',
	'≸',
	'&ntlg;',
	'⋪',
	'&ntriangleleft;',
	'⋬',
	'&ntrianglelefteq;',
	'⋫',
	'&ntriangleright;',
	'⋭',
	'&ntrianglerighteq;',
	'Ν',
	'&Nu;',
	'ν',
	'&nu;',
	'#',
	'&num;',
	'№',
	'&numero;',
	' ',
	'&numsp;',
	'≍⃒',
	'&nvap;',
	'⊯',
	'&nVDash;',
	'⊮',
	'&nVdash;',
	'⊭',
	'&nvDash;',
	'⊬',
	'&nvdash;',
	'≥⃒',
	'&nvge;',
	'>⃒',
	'&nvgt;',
	'⤄',
	'&nvHarr;',
	'⧞',
	'&nvinfin;',
	'⤂',
	'&nvlArr;',
	'≤⃒',
	'&nvle;',
	'<⃒',
	'&nvlt;',
	'⊴⃒',
	'&nvltrie;',
	'⤃',
	'&nvrArr;',
	'⊵⃒',
	'&nvrtrie;',
	'∼⃒',
	'&nvsim;',
	'⤣',
	'&nwarhk;',
	'⇖',
	'&nwArr;',
	'↖',
	'&nwarr;',
	'↖',
	'&nwarrow;',
	'⤧',
	'&nwnear;',
	'Ó',
	'&Oacute;',
	'ó',
	'&oacute;',
	'⊛',
	'&oast;',
	'⊚',
	'&ocir;',
	'Ô',
	'&Ocirc;',
	'ô',
	'&ocirc;',
	'О',
	'&Ocy;',
	'о',
	'&ocy;',
	'⊝',
	'&odash;',
	'Ő',
	'&Odblac;',
	'ő',
	'&odblac;',
	'⨸',
	'&odiv;',
	'⊙',
	'&odot;',
	'⦼',
	'&odsold;',
	'Œ',
	'&OElig;',
	'œ',
	'&oelig;',
	'⦿',
	'&ofcir;',
	'𝔒',
	'&Ofr;',
	'𝔬',
	'&ofr;',
	'˛',
	'&ogon;',
	'Ò',
	'&Ograve;',
	'ò',
	'&ograve;',
	'⧁',
	'&ogt;',
	'⦵',
	'&ohbar;',
	'Ω',
	'&ohm;',
	'∮',
	'&oint;',
	'↺',
	'&olarr;',
	'⦾',
	'&olcir;',
	'⦻',
	'&olcross;',
	'‾',
	'&oline;',
	'⧀',
	'&olt;',
	'Ō',
	'&Omacr;',
	'ō',
	'&omacr;',
	'Ω',
	'&Omega;',
	'ω',
	'&omega;',
	'Ο',
	'&Omicron;',
	'ο',
	'&omicron;',
	'⦶',
	'&omid;',
	'⊖',
	'&ominus;',
	'𝕆',
	'&Oopf;',
	'𝕠',
	'&oopf;',
	'⦷',
	'&opar;',
	'“',
	'&OpenCurlyDoubleQuote;',
	'‘',
	'&OpenCurlyQuote;',
	'⦹',
	'&operp;',
	'⊕',
	'&oplus;',
	'⩔',
	'&Or;',
	'∨',
	'&or;',
	'↻',
	'&orarr;',
	'⩝',
	'&ord;',
	'ℴ',
	'&order;',
	'ℴ',
	'&orderof;',
	'ª',
	'&ordf;',
	'º',
	'&ordm;',
	'⊶',
	'&origof;',
	'⩖',
	'&oror;',
	'⩗',
	'&orslope;',
	'⩛',
	'&orv;',
	'Ⓢ',
	'&oS;',
	'𝒪',
	'&Oscr;',
	'ℴ',
	'&oscr;',
	'Ø',
	'&Oslash;',
	'ø',
	'&oslash;',
	'⊘',
	'&osol;',
	'Õ',
	'&Otilde;',
	'õ',
	'&otilde;',
	'⨷',
	'&Otimes;',
	'⊗',
	'&otimes;',
	'⨶',
	'&otimesas;',
	'Ö',
	'&Ouml;',
	'ö',
	'&ouml;',
	'⌽',
	'&ovbar;',
	'‾',
	'&OverBar;',
	'⏞',
	'&OverBrace;',
	'⎴',
	'&OverBracket;',
	'⏜',
	'&OverParenthesis;',
	'∥',
	'&par;',
	'¶',
	'&para;',
	'∥',
	'&parallel;',
	'⫳',
	'&parsim;',
	'⫽',
	'&parsl;',
	'∂',
	'&part;',
	'∂',
	'&PartialD;',
	'П',
	'&Pcy;',
	'п',
	'&pcy;',
	'%',
	'&percnt;',
	'.',
	'&period;',
	'‰',
	'&permil;',
	'⊥',
	'&perp;',
	'‱',
	'&pertenk;',
	'𝔓',
	'&Pfr;',
	'𝔭',
	'&pfr;',
	'Φ',
	'&Phi;',
	'φ',
	'&phi;',
	'ϕ',
	'&phiv;',
	'ℳ',
	'&phmmat;',
	'☎',
	'&phone;',
	'Π',
	'&Pi;',
	'π',
	'&pi;',
	'⋔',
	'&pitchfork;',
	'ϖ',
	'&piv;',
	'ℏ',
	'&planck;',
	'ℎ',
	'&planckh;',
	'ℏ',
	'&plankv;',
	'+',
	'&plus;',
	'⨣',
	'&plusacir;',
	'⊞',
	'&plusb;',
	'⨢',
	'&pluscir;',
	'∔',
	'&plusdo;',
	'⨥',
	'&plusdu;',
	'⩲',
	'&pluse;',
	'±',
	'&PlusMinus;',
	'±',
	'&plusmn;',
	'⨦',
	'&plussim;',
	'⨧',
	'&plustwo;',
	'±',
	'&pm;',
	'ℌ',
	'&Poincareplane;',
	'⨕',
	'&pointint;',
	'ℙ',
	'&Popf;',
	'𝕡',
	'&popf;',
	'£',
	'&pound;',
	'⪻',
	'&Pr;',
	'≺',
	'&pr;',
	'⪷',
	'&prap;',
	'≼',
	'&prcue;',
	'⪳',
	'&prE;',
	'⪯',
	'&pre;',
	'≺',
	'&prec;',
	'⪷',
	'&precapprox;',
	'≼',
	'&preccurlyeq;',
	'≺',
	'&Precedes;',
	'⪯',
	'&PrecedesEqual;',
	'≼',
	'&PrecedesSlantEqual;',
	'≾',
	'&PrecedesTilde;',
	'⪯',
	'&preceq;',
	'⪹',
	'&precnapprox;',
	'⪵',
	'&precneqq;',
	'⋨',
	'&precnsim;',
	'≾',
	'&precsim;',
	'″',
	'&Prime;',
	'′',
	'&prime;',
	'ℙ',
	'&primes;',
	'⪹',
	'&prnap;',
	'⪵',
	'&prnE;',
	'⋨',
	'&prnsim;',
	'∏',
	'&prod;',
	'∏',
	'&Product;',
	'⌮',
	'&profalar;',
	'⌒',
	'&profline;',
	'⌓',
	'&profsurf;',
	'∝',
	'&prop;',
	'∷',
	'&Proportion;',
	'∝',
	'&Proportional;',
	'∝',
	'&propto;',
	'≾',
	'&prsim;',
	'⊰',
	'&prurel;',
	'𝒫',
	'&Pscr;',
	'𝓅',
	'&pscr;',
	'Ψ',
	'&Psi;',
	'ψ',
	'&psi;',
	' ',
	'&puncsp;',
	'𝔔',
	'&Qfr;',
	'𝔮',
	'&qfr;',
	'⨌',
	'&qint;',
	'ℚ',
	'&Qopf;',
	'𝕢',
	'&qopf;',
	'⁗',
	'&qprime;',
	'𝒬',
	'&Qscr;',
	'𝓆',
	'&qscr;',
	'ℍ',
	'&quaternions;',
	'⨖',
	'&quatint;',
	'?',
	'&quest;',
	'≟',
	'&questeq;',
	'"',
	'&QUOT;',
	'"',
	'&quot;',
	'⇛',
	'&rAarr;',
	'∽̱',
	'&race;',
	'Ŕ',
	'&Racute;',
	'ŕ',
	'&racute;',
	'√',
	'&radic;',
	'⦳',
	'&raemptyv;',
	'⟫',
	'&Rang;',
	'⟩',
	'&rang;',
	'⦒',
	'&rangd;',
	'⦥',
	'&range;',
	'⟩',
	'&rangle;',
	'»',
	'&raquo;',
	'↠',
	'&Rarr;',
	'⇒',
	'&rArr;',
	'→',
	'&rarr;',
	'⥵',
	'&rarrap;',
	'⇥',
	'&rarrb;',
	'⤠',
	'&rarrbfs;',
	'⤳',
	'&rarrc;',
	'⤞',
	'&rarrfs;',
	'↪',
	'&rarrhk;',
	'↬',
	'&rarrlp;',
	'⥅',
	'&rarrpl;',
	'⥴',
	'&rarrsim;',
	'⤖',
	'&Rarrtl;',
	'↣',
	'&rarrtl;',
	'↝',
	'&rarrw;',
	'⤜',
	'&rAtail;',
	'⤚',
	'&ratail;',
	'∶',
	'&ratio;',
	'ℚ',
	'&rationals;',
	'⤐',
	'&RBarr;',
	'⤏',
	'&rBarr;',
	'⤍',
	'&rbarr;',
	'❳',
	'&rbbrk;',
	'}',
	'&rbrace;',
	']',
	'&rbrack;',
	'⦌',
	'&rbrke;',
	'⦎',
	'&rbrksld;',
	'⦐',
	'&rbrkslu;',
	'Ř',
	'&Rcaron;',
	'ř',
	'&rcaron;',
	'Ŗ',
	'&Rcedil;',
	'ŗ',
	'&rcedil;',
	'⌉',
	'&rceil;',
	'}',
	'&rcub;',
	'Р',
	'&Rcy;',
	'р',
	'&rcy;',
	'⤷',
	'&rdca;',
	'⥩',
	'&rdldhar;',
	'”',
	'&rdquo;',
	'”',
	'&rdquor;',
	'↳',
	'&rdsh;',
	'ℜ',
	'&Re;',
	'ℜ',
	'&real;',
	'ℛ',
	'&realine;',
	'ℜ',
	'&realpart;',
	'ℝ',
	'&reals;',
	'▭',
	'&rect;',
	'®',
	'&REG;',
	'®',
	'&reg;',
	'∋',
	'&ReverseElement;',
	'⇋',
	'&ReverseEquilibrium;',
	'⥯',
	'&ReverseUpEquilibrium;',
	'⥽',
	'&rfisht;',
	'⌋',
	'&rfloor;',
	'ℜ',
	'&Rfr;',
	'𝔯',
	'&rfr;',
	'⥤',
	'&rHar;',
	'⇁',
	'&rhard;',
	'⇀',
	'&rharu;',
	'⥬',
	'&rharul;',
	'Ρ',
	'&Rho;',
	'ρ',
	'&rho;',
	'ϱ',
	'&rhov;',
	'⟩',
	'&RightAngleBracket;',
	'→',
	'&RightArrow;',
	'⇒',
	'&Rightarrow;',
	'→',
	'&rightarrow;',
	'⇥',
	'&RightArrowBar;',
	'⇄',
	'&RightArrowLeftArrow;',
	'↣',
	'&rightarrowtail;',
	'⌉',
	'&RightCeiling;',
	'⟧',
	'&RightDoubleBracket;',
	'⥝',
	'&RightDownTeeVector;',
	'⇂',
	'&RightDownVector;',
	'⥕',
	'&RightDownVectorBar;',
	'⌋',
	'&RightFloor;',
	'⇁',
	'&rightharpoondown;',
	'⇀',
	'&rightharpoonup;',
	'⇄',
	'&rightleftarrows;',
	'⇌',
	'&rightleftharpoons;',
	'⇉',
	'&rightrightarrows;',
	'↝',
	'&rightsquigarrow;',
	'⊢',
	'&RightTee;',
	'↦',
	'&RightTeeArrow;',
	'⥛',
	'&RightTeeVector;',
	'⋌',
	'&rightthreetimes;',
	'⊳',
	'&RightTriangle;',
	'⧐',
	'&RightTriangleBar;',
	'⊵',
	'&RightTriangleEqual;',
	'⥏',
	'&RightUpDownVector;',
	'⥜',
	'&RightUpTeeVector;',
	'↾',
	'&RightUpVector;',
	'⥔',
	'&RightUpVectorBar;',
	'⇀',
	'&RightVector;',
	'⥓',
	'&RightVectorBar;',
	'˚',
	'&ring;',
	'≓',
	'&risingdotseq;',
	'⇄',
	'&rlarr;',
	'⇌',
	'&rlhar;',
	'‏',
	'&rlm;',
	'⎱',
	'&rmoust;',
	'⎱',
	'&rmoustache;',
	'⫮',
	'&rnmid;',
	'⟭',
	'&roang;',
	'⇾',
	'&roarr;',
	'⟧',
	'&robrk;',
	'⦆',
	'&ropar;',
	'ℝ',
	'&Ropf;',
	'𝕣',
	'&ropf;',
	'⨮',
	'&roplus;',
	'⨵',
	'&rotimes;',
	'⥰',
	'&RoundImplies;',
	')',
	'&rpar;',
	'⦔',
	'&rpargt;',
	'⨒',
	'&rppolint;',
	'⇉',
	'&rrarr;',
	'⇛',
	'&Rrightarrow;',
	'›',
	'&rsaquo;',
	'ℛ',
	'&Rscr;',
	'𝓇',
	'&rscr;',
	'↱',
	'&Rsh;',
	'↱',
	'&rsh;',
	']',
	'&rsqb;',
	'’',
	'&rsquo;',
	'’',
	'&rsquor;',
	'⋌',
	'&rthree;',
	'⋊',
	'&rtimes;',
	'▹',
	'&rtri;',
	'⊵',
	'&rtrie;',
	'▸',
	'&rtrif;',
	'⧎',
	'&rtriltri;',
	'⧴',
	'&RuleDelayed;',
	'⥨',
	'&ruluhar;',
	'℞',
	'&rx;',
	'Ś',
	'&Sacute;',
	'ś',
	'&sacute;',
	'‚',
	'&sbquo;',
	'⪼',
	'&Sc;',
	'≻',
	'&sc;',
	'⪸',
	'&scap;',
	'Š',
	'&Scaron;',
	'š',
	'&scaron;',
	'≽',
	'&sccue;',
	'⪴',
	'&scE;',
	'⪰',
	'&sce;',
	'Ş',
	'&Scedil;',
	'ş',
	'&scedil;',
	'Ŝ',
	'&Scirc;',
	'ŝ',
	'&scirc;',
	'⪺',
	'&scnap;',
	'⪶',
	'&scnE;',
	'⋩',
	'&scnsim;',
	'⨓',
	'&scpolint;',
	'≿',
	'&scsim;',
	'С',
	'&Scy;',
	'с',
	'&scy;',
	'⋅',
	'&sdot;',
	'⊡',
	'&sdotb;',
	'⩦',
	'&sdote;',
	'⤥',
	'&searhk;',
	'⇘',
	'&seArr;',
	'↘',
	'&searr;',
	'↘',
	'&searrow;',
	'§',
	'&sect;',
	';',
	'&semi;',
	'⤩',
	'&seswar;',
	'∖',
	'&setminus;',
	'∖',
	'&setmn;',
	'✶',
	'&sext;',
	'𝔖',
	'&Sfr;',
	'𝔰',
	'&sfr;',
	'⌢',
	'&sfrown;',
	'♯',
	'&sharp;',
	'Щ',
	'&SHCHcy;',
	'щ',
	'&shchcy;',
	'Ш',
	'&SHcy;',
	'ш',
	'&shcy;',
	'↓',
	'&ShortDownArrow;',
	'←',
	'&ShortLeftArrow;',
	'∣',
	'&shortmid;',
	'∥',
	'&shortparallel;',
	'→',
	'&ShortRightArrow;',
	'↑',
	'&ShortUpArrow;',
	'­',
	'&shy;',
	'Σ',
	'&Sigma;',
	'σ',
	'&sigma;',
	'ς',
	'&sigmaf;',
	'ς',
	'&sigmav;',
	'∼',
	'&sim;',
	'⩪',
	'&simdot;',
	'≃',
	'&sime;',
	'≃',
	'&simeq;',
	'⪞',
	'&simg;',
	'⪠',
	'&simgE;',
	'⪝',
	'&siml;',
	'⪟',
	'&simlE;',
	'≆',
	'&simne;',
	'⨤',
	'&simplus;',
	'⥲',
	'&simrarr;',
	'←',
	'&slarr;',
	'∘',
	'&SmallCircle;',
	'∖',
	'&smallsetminus;',
	'⨳',
	'&smashp;',
	'⧤',
	'&smeparsl;',
	'∣',
	'&smid;',
	'⌣',
	'&smile;',
	'⪪',
	'&smt;',
	'⪬',
	'&smte;',
	'⪬︀',
	'&smtes;',
	'Ь',
	'&SOFTcy;',
	'ь',
	'&softcy;',
	'/',
	'&sol;',
	'⧄',
	'&solb;',
	'⌿',
	'&solbar;',
	'𝕊',
	'&Sopf;',
	'𝕤',
	'&sopf;',
	'♠',
	'&spades;',
	'♠',
	'&spadesuit;',
	'∥',
	'&spar;',
	'⊓',
	'&sqcap;',
	'⊓︀',
	'&sqcaps;',
	'⊔',
	'&sqcup;',
	'⊔︀',
	'&sqcups;',
	'√',
	'&Sqrt;',
	'⊏',
	'&sqsub;',
	'⊑',
	'&sqsube;',
	'⊏',
	'&sqsubset;',
	'⊑',
	'&sqsubseteq;',
	'⊐',
	'&sqsup;',
	'⊒',
	'&sqsupe;',
	'⊐',
	'&sqsupset;',
	'⊒',
	'&sqsupseteq;',
	'□',
	'&squ;',
	'□',
	'&Square;',
	'□',
	'&square;',
	'⊓',
	'&SquareIntersection;',
	'⊏',
	'&SquareSubset;',
	'⊑',
	'&SquareSubsetEqual;',
	'⊐',
	'&SquareSuperset;',
	'⊒',
	'&SquareSupersetEqual;',
	'⊔',
	'&SquareUnion;',
	'▪',
	'&squarf;',
	'▪',
	'&squf;',
	'→',
	'&srarr;',
	'𝒮',
	'&Sscr;',
	'𝓈',
	'&sscr;',
	'∖',
	'&ssetmn;',
	'⌣',
	'&ssmile;',
	'⋆',
	'&sstarf;',
	'⋆',
	'&Star;',
	'☆',
	'&star;',
	'★',
	'&starf;',
	'ϵ',
	'&straightepsilon;',
	'ϕ',
	'&straightphi;',
	'¯',
	'&strns;',
	'⋐',
	'&Sub;',
	'⊂',
	'&sub;',
	'⪽',
	'&subdot;',
	'⫅',
	'&subE;',
	'⊆',
	'&sube;',
	'⫃',
	'&subedot;',
	'⫁',
	'&submult;',
	'⫋',
	'&subnE;',
	'⊊',
	'&subne;',
	'⪿',
	'&subplus;',
	'⥹',
	'&subrarr;',
	'⋐',
	'&Subset;',
	'⊂',
	'&subset;',
	'⊆',
	'&subseteq;',
	'⫅',
	'&subseteqq;',
	'⊆',
	'&SubsetEqual;',
	'⊊',
	'&subsetneq;',
	'⫋',
	'&subsetneqq;',
	'⫇',
	'&subsim;',
	'⫕',
	'&subsub;',
	'⫓',
	'&subsup;',
	'≻',
	'&succ;',
	'⪸',
	'&succapprox;',
	'≽',
	'&succcurlyeq;',
	'≻',
	'&Succeeds;',
	'⪰',
	'&SucceedsEqual;',
	'≽',
	'&SucceedsSlantEqual;',
	'≿',
	'&SucceedsTilde;',
	'⪰',
	'&succeq;',
	'⪺',
	'&succnapprox;',
	'⪶',
	'&succneqq;',
	'⋩',
	'&succnsim;',
	'≿',
	'&succsim;',
	'∋',
	'&SuchThat;',
	'∑',
	'&Sum;',
	'∑',
	'&sum;',
	'♪',
	'&sung;',
	'⋑',
	'&Sup;',
	'⊃',
	'&sup;',
	'¹',
	'&sup1;',
	'²',
	'&sup2;',
	'³',
	'&sup3;',
	'⪾',
	'&supdot;',
	'⫘',
	'&supdsub;',
	'⫆',
	'&supE;',
	'⊇',
	'&supe;',
	'⫄',
	'&supedot;',
	'⊃',
	'&Superset;',
	'⊇',
	'&SupersetEqual;',
	'⟉',
	'&suphsol;',
	'⫗',
	'&suphsub;',
	'⥻',
	'&suplarr;',
	'⫂',
	'&supmult;',
	'⫌',
	'&supnE;',
	'⊋',
	'&supne;',
	'⫀',
	'&supplus;',
	'⋑',
	'&Supset;',
	'⊃',
	'&supset;',
	'⊇',
	'&supseteq;',
	'⫆',
	'&supseteqq;',
	'⊋',
	'&supsetneq;',
	'⫌',
	'&supsetneqq;',
	'⫈',
	'&supsim;',
	'⫔',
	'&supsub;',
	'⫖',
	'&supsup;',
	'⤦',
	'&swarhk;',
	'⇙',
	'&swArr;',
	'↙',
	'&swarr;',
	'↙',
	'&swarrow;',
	'⤪',
	'&swnwar;',
	'ß',
	'&szlig;',
	'␉',
	'&Tab;',
	'⌖',
	'&target;',
	'Τ',
	'&Tau;',
	'τ',
	'&tau;',
	'⎴',
	'&tbrk;',
	'Ť',
	'&Tcaron;',
	'ť',
	'&tcaron;',
	'Ţ',
	'&Tcedil;',
	'ţ',
	'&tcedil;',
	'Т',
	'&Tcy;',
	'т',
	'&tcy;',
	'◌⃛',
	'&tdot;',
	'⌕',
	'&telrec;',
	'𝔗',
	'&Tfr;',
	'𝔱',
	'&tfr;',
	'∴',
	'&there4;',
	'∴',
	'&Therefore;',
	'∴',
	'&therefore;',
	'Θ',
	'&Theta;',
	'θ',
	'&theta;',
	'ϑ',
	'&thetasym;',
	'ϑ',
	'&thetav;',
	'≈',
	'&thickapprox;',
	'∼',
	'&thicksim;',
	'  ',
	'&ThickSpace;',
	' ',
	'&thinsp;',
	' ',
	'&ThinSpace;',
	'≈',
	'&thkap;',
	'∼',
	'&thksim;',
	'Þ',
	'&THORN;',
	'þ',
	'&thorn;',
	'∼',
	'&Tilde;',
	'˜',
	'&tilde;',
	'≃',
	'&TildeEqual;',
	'≅',
	'&TildeFullEqual;',
	'≈',
	'&TildeTilde;',
	'×',
	'&times;',
	'⊠',
	'&timesb;',
	'⨱',
	'&timesbar;',
	'⨰',
	'&timesd;',
	'∭',
	'&tint;',
	'⤨',
	'&toea;',
	'⊤',
	'&top;',
	'⌶',
	'&topbot;',
	'⫱',
	'&topcir;',
	'𝕋',
	'&Topf;',
	'𝕥',
	'&topf;',
	'⫚',
	'&topfork;',
	'⤩',
	'&tosa;',
	'‴',
	'&tprime;',
	'™',
	'&TRADE;',
	'™',
	'&trade;',
	'▵',
	'&triangle;',
	'▿',
	'&triangledown;',
	'◃',
	'&triangleleft;',
	'⊴',
	'&trianglelefteq;',
	'≜',
	'&triangleq;',
	'▹',
	'&triangleright;',
	'⊵',
	'&trianglerighteq;',
	'◬',
	'&tridot;',
	'≜',
	'&trie;',
	'⨺',
	'&triminus;',
	'◌⃛',
	'&TripleDot;',
	'⨹',
	'&triplus;',
	'⧍',
	'&trisb;',
	'⨻',
	'&tritime;',
	'⏢',
	'&trpezium;',
	'𝒯',
	'&Tscr;',
	'𝓉',
	'&tscr;',
	'Ц',
	'&TScy;',
	'ц',
	'&tscy;',
	'Ћ',
	'&TSHcy;',
	'ћ',
	'&tshcy;',
	'Ŧ',
	'&Tstrok;',
	'ŧ',
	'&tstrok;',
	'≬',
	'&twixt;',
	'↞',
	'&twoheadleftarrow;',
	'↠',
	'&twoheadrightarrow;',
	'Ú',
	'&Uacute;',
	'ú',
	'&uacute;',
	'↟',
	'&Uarr;',
	'⇑',
	'&uArr;',
	'↑',
	'&uarr;',
	'⥉',
	'&Uarrocir;',
	'Ў',
	'&Ubrcy;',
	'ў',
	'&ubrcy;',
	'Ŭ',
	'&Ubreve;',
	'ŭ',
	'&ubreve;',
	'Û',
	'&Ucirc;',
	'û',
	'&ucirc;',
	'У',
	'&Ucy;',
	'у',
	'&ucy;',
	'⇅',
	'&udarr;',
	'Ű',
	'&Udblac;',
	'ű',
	'&udblac;',
	'⥮',
	'&udhar;',
	'⥾',
	'&ufisht;',
	'𝔘',
	'&Ufr;',
	'𝔲',
	'&ufr;',
	'Ù',
	'&Ugrave;',
	'ù',
	'&ugrave;',
	'⥣',
	'&uHar;',
	'↿',
	'&uharl;',
	'↾',
	'&uharr;',
	'▀',
	'&uhblk;',
	'⌜',
	'&ulcorn;',
	'⌜',
	'&ulcorner;',
	'⌏',
	'&ulcrop;',
	'◸',
	'&ultri;',
	'Ū',
	'&Umacr;',
	'ū',
	'&umacr;',
	'¨',
	'&uml;',
	'_',
	'&UnderBar;',
	'⏟',
	'&UnderBrace;',
	'⎵',
	'&UnderBracket;',
	'⏝',
	'&UnderParenthesis;',
	'⋃',
	'&Union;',
	'⊎',
	'&UnionPlus;',
	'Ų',
	'&Uogon;',
	'ų',
	'&uogon;',
	'𝕌',
	'&Uopf;',
	'𝕦',
	'&uopf;',
	'↑',
	'&UpArrow;',
	'⇑',
	'&Uparrow;',
	'↑',
	'&uparrow;',
	'⤒',
	'&UpArrowBar;',
	'⇅',
	'&UpArrowDownArrow;',
	'↕',
	'&UpDownArrow;',
	'⇕',
	'&Updownarrow;',
	'↕',
	'&updownarrow;',
	'⥮',
	'&UpEquilibrium;',
	'↿',
	'&upharpoonleft;',
	'↾',
	'&upharpoonright;',
	'⊎',
	'&uplus;',
	'↖',
	'&UpperLeftArrow;',
	'↗',
	'&UpperRightArrow;',
	'ϒ',
	'&Upsi;',
	'υ',
	'&upsi;',
	'ϒ',
	'&upsih;',
	'Υ',
	'&Upsilon;',
	'υ',
	'&upsilon;',
	'⊥',
	'&UpTee;',
	'↥',
	'&UpTeeArrow;',
	'⇈',
	'&upuparrows;',
	'⌝',
	'&urcorn;',
	'⌝',
	'&urcorner;',
	'⌎',
	'&urcrop;',
	'Ů',
	'&Uring;',
	'ů',
	'&uring;',
	'◹',
	'&urtri;',
	'𝒰',
	'&Uscr;',
	'𝓊',
	'&uscr;',
	'⋰',
	'&utdot;',
	'Ũ',
	'&Utilde;',
	'ũ',
	'&utilde;',
	'▵',
	'&utri;',
	'▴',
	'&utrif;',
	'⇈',
	'&uuarr;',
	'Ü',
	'&Uuml;',
	'ü',
	'&uuml;',
	'⦧',
	'&uwangle;',
	'⦜',
	'&vangrt;',
	'ϵ',
	'&varepsilon;',
	'ϰ',
	'&varkappa;',
	'∅',
	'&varnothing;',
	'ϕ',
	'&varphi;',
	'ϖ',
	'&varpi;',
	'∝',
	'&varpropto;',
	'⇕',
	'&vArr;',
	'↕',
	'&varr;',
	'ϱ',
	'&varrho;',
	'ς',
	'&varsigma;',
	'⊊︀',
	'&varsubsetneq;',
	'⫋︀',
	'&varsubsetneqq;',
	'⊋︀',
	'&varsupsetneq;',
	'⫌︀',
	'&varsupsetneqq;',
	'ϑ',
	'&vartheta;',
	'⊲',
	'&vartriangleleft;',
	'⊳',
	'&vartriangleright;',
	'⫫',
	'&Vbar;',
	'⫨',
	'&vBar;',
	'⫩',
	'&vBarv;',
	'В',
	'&Vcy;',
	'в',
	'&vcy;',
	'⊫',
	'&VDash;',
	'⊩',
	'&Vdash;',
	'⊨',
	'&vDash;',
	'⊢',
	'&vdash;',
	'⫦',
	'&Vdashl;',
	'⋁',
	'&Vee;',
	'∨',
	'&vee;',
	'⊻',
	'&veebar;',
	'≚',
	'&veeeq;',
	'⋮',
	'&vellip;',
	'‖',
	'&Verbar;',
	'|',
	'&verbar;',
	'‖',
	'&Vert;',
	'|',
	'&vert;',
	'∣',
	'&VerticalBar;',
	'|',
	'&VerticalLine;',
	'❘',
	'&VerticalSeparator;',
	'≀',
	'&VerticalTilde;',
	' ',
	'&VeryThinSpace;',
	'𝔙',
	'&Vfr;',
	'𝔳',
	'&vfr;',
	'⊲',
	'&vltri;',
	'⊂⃒',
	'&vnsub;',
	'⊃⃒',
	'&vnsup;',
	'𝕍',
	'&Vopf;',
	'𝕧',
	'&vopf;',
	'∝',
	'&vprop;',
	'⊳',
	'&vrtri;',
	'𝒱',
	'&Vscr;',
	'𝓋',
	'&vscr;',
	'⫋︀',
	'&vsubnE;',
	'⊊︀',
	'&vsubne;',
	'⫌︀',
	'&vsupnE;',
	'⊋︀',
	'&vsupne;',
	'⊪',
	'&Vvdash;',
	'⦚',
	'&vzigzag;',
	'Ŵ',
	'&Wcirc;',
	'ŵ',
	'&wcirc;',
	'⩟',
	'&wedbar;',
	'⋀',
	'&Wedge;',
	'∧',
	'&wedge;',
	'≙',
	'&wedgeq;',
	'℘',
	'&weierp;',
	'𝔚',
	'&Wfr;',
	'𝔴',
	'&wfr;',
	'𝕎',
	'&Wopf;',
	'𝕨',
	'&wopf;',
	'℘',
	'&wp;',
	'≀',
	'&wr;',
	'≀',
	'&wreath;',
	'𝒲',
	'&Wscr;',
	'𝓌',
	'&wscr;',
	'⋂',
	'&xcap;',
	'◯',
	'&xcirc;',
	'⋃',
	'&xcup;',
	'▽',
	'&xdtri;',
	'𝔛',
	'&Xfr;',
	'𝔵',
	'&xfr;',
	'⟺',
	'&xhArr;',
	'⟷',
	'&xharr;',
	'Ξ',
	'&Xi;',
	'ξ',
	'&xi;',
	'⟸',
	'&xlArr;',
	'⟵',
	'&xlarr;',
	'⟼',
	'&xmap;',
	'⋻',
	'&xnis;',
	'⨀',
	'&xodot;',
	'𝕏',
	'&Xopf;',
	'𝕩',
	'&xopf;',
	'⨁',
	'&xoplus;',
	'⨂',
	'&xotime;',
	'⟹',
	'&xrArr;',
	'⟶',
	'&xrarr;',
	'𝒳',
	'&Xscr;',
	'𝓍',
	'&xscr;',
	'⨆',
	'&xsqcup;',
	'⨄',
	'&xuplus;',
	'△',
	'&xutri;',
	'⋁',
	'&xvee;',
	'⋀',
	'&xwedge;',
	'Ý',
	'&Yacute;',
	'ý',
	'&yacute;',
	'Я',
	'&YAcy;',
	'я',
	'&yacy;',
	'Ŷ',
	'&Ycirc;',
	'ŷ',
	'&ycirc;',
	'Ы',
	'&Ycy;',
	'ы',
	'&ycy;',
	'¥',
	'&yen;',
	'𝔜',
	'&Yfr;',
	'𝔶',
	'&yfr;',
	'Ї',
	'&YIcy;',
	'ї',
	'&yicy;',
	'𝕐',
	'&Yopf;',
	'𝕪',
	'&yopf;',
	'𝒴',
	'&Yscr;',
	'𝓎',
	'&yscr;',
	'Ю',
	'&YUcy;',
	'ю',
	'&yucy;',
	'Ÿ',
	'&Yuml;',
	'ÿ',
	'&yuml;',
	'Ź',
	'&Zacute;',
	'ź',
	'&zacute;',
	'Ž',
	'&Zcaron;',
	'ž',
	'&zcaron;',
	'З',
	'&Zcy;',
	'з',
	'&zcy;',
	'Ż',
	'&Zdot;',
	'ż',
	'&zdot;',
	'ℨ',
	'&zeetrf;',
	'​',
	'&ZeroWidthSpace;',
	'Ζ',
	'&Zeta;',
	'ζ',
	'&zeta;',
	'ℨ',
	'&Zfr;',
	'𝔷',
	'&zfr;',
	'Ж',
	'&ZHcy;',
	'ж',
	'&zhcy;',
	'⇝',
	'&zigrarr;',
	'ℤ',
	'&Zopf;',
	'𝕫',
	'&zopf;',
	'𝒵',
	'&Zscr;',
	'𝓏',
	'&zscr;',
	'‍',
	'&zwj;',
	'‌',
	'&zwnj;',
]
